

module dc(clk, en, x, y);
input clk, en;
input [23:0] x;
output reg [7:0] y;

wire sys_clk = clk;
wire sys_en = en;

always @(posedge sys_clk, negedge sys_en) begin
if(~sys_en)begin
	y = 8'b0;
end else begin

case(x) 
24'b	0101110	:	y=	8'h41	;
24'b	01110101010	:	y=	8'h42	;
24'b	0111010111010	:	y=	8'h43	;
24'b	011101010	:	y=	8'h44	;
24'b	010	:	y=	8'h45	;
24'b	01010111010	:	y=	8'h46	;
24'b	01110111010	:	y=	8'h47	;
24'b	010101010	:	y=	8'h48	;
24'b	01010	:	y=	8'h49	;
24'b	010111011101110	:	y=	8'h4A	;
24'b	01110101110	:	y=	8'h4B	;
24'b	0101110101	:	y=	8'h4C	;
24'b	011101110	:	y=	8'h4D	;
24'b	0111010	:	y=	8'h4E	;
24'b	0111011101110	:	y=	8'h4F	;
24'b	010111011101	:	y=	8'h50	;
24'b	011101110101110	:	y=	8'h51	;
24'b	010111010	:	y=	8'h52	;
24'b	0101010	:	y=	8'h53	;
24'b	01110	:	y=	8'h54	;
24'b	010101110	:	y=	8'h55	;
24'b	01010101110	:	y=	8'h56	;
24'b	01011101110	:	y=	8'h57	;
24'b	0111010101110	:	y=	8'h58	;
24'b	011101011101110	:	y=	8'h59	;
24'b	0111011101010	:	y=	8'h5A	;
					
					
24'b	0101110111011101110	:	y=	8'h31	;
24'b	01010111011101110	:	y=	8'h32	;
24'b	010101011101110	:	y=	8'h33	;
24'b	0101010101110	:	y=	8'h34	;
24'b	01010101010	:	y=	8'h35	;
24'b	0111010101010	:	y=	8'h36	;
24'b	011101110101010	:	y=	8'h37	;
24'b	01110111011101010	:	y=	8'h38	;
24'b	0111011101110111010	:	y=	8'h39	;
24'b	011101110111011101110	:	y=	8'h30	;
24'b	0101010101010	:	y=	8'h2E	;
24'b	0101110101110101110	:	y=	8'h2C	;
24'b	011101110111010101	:	y=	8'h3A	;
24'b	0111010111010111010	:	y=	8'h3B	;
24'b	011101011101110101110	:	y=	8'h28	;
24'b	010111011101110111010	:	y=	8'h27	;
24'b	01011101010111010	:	y=	8'h22	;
24'b	01110101010101110	:	y=	8'h2D	;
24'b	011101010111010	:	y=	8'h2F	;
24'b	0101011101110101110	:	y=	8'h5F	;
24'b	0101011101110101	:	y=	8'h3F	;
24'b	01110111010101110111	:	y=	8'h21	;
24'b	010111010111010	:	y=	8'h2B	;

24'b	0101110111010111010	:	y=	8'h40	;
24'b	010101110101110	:	y=	8'hFF	;
24'b	0	:	y=	8'h20	;


default y=8'b0;

endcase

end

end

endmodule
